// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this
// file, You can obtain one at http://mozilla.org/MPL/2.0/.

module cc
import gg

pub struct BaseApp {
}

fn (mut app BaseApp) setup() {}
fn (mut app BaseApp) update() {}
fn (mut app BaseApp) draw() {}
fn (mut app BaseApp) on_event(event &gg.Event) {}
fn (mut app BaseApp) key_pressed(keycode gg.KeyCode, m gg.Modifier) {}
fn (mut app BaseApp) key_released(keycode gg.KeyCode, m gg.Modifier) {}
fn (mut app BaseApp) mouse_pressed(x f32, y f32, button gg.MouseButton) {}
fn (mut app BaseApp) mouse_released(x f32, y f32, button gg.MouseButton) {}
fn (mut app BaseApp) mouse_moved(x f32, y f32) {}
fn (mut app BaseApp) exit() {}

interface IApp {
mut:
	setup()
	update()
	draw()
	on_event(&gg.Event)
	key_pressed(gg.KeyCode, gg.Modifier)
	key_released(gg.KeyCode, gg.Modifier)
	mouse_pressed(f32, f32, gg.MouseButton)
	mouse_released(f32, f32, gg.MouseButton)
	mouse_moved(f32, f32)
	exit()
}
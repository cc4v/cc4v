// Reference:
// https://github.com/openframeworks/openFrameworks/blob/996f7880bc250254480561a2f2dab3554a830084/libs/openFrameworks/gl/ofGLProgrammableRenderer.cpp

module cc
// import gg
import sokol.sgl
import log

const cc_max_style_history = 32

pub fn push_matrix() {
	sgl.push_matrix()
}

pub fn pop_matrix() {
	sgl.pop_matrix()
}

fn set_style(style &CCStyle, mut c CC) {
	c.current_style = style
}

pub fn push_style() {
	sgl.push_pipeline()

	mut ctx := context()
	if unsafe { ctx.cc == nil } {
		ctx.cc.style_history.push(ctx.cc.current_style)
		if ctx.cc.style_history.len() > cc_max_style_history {
			ctx.cc.style_history.pop() or { panic(err) }
			log.warn("cc: push_style() maximum number of style pushes ${cc_max_style_history} reached, did you forget to pop somewhere?")
		}
	}
}

pub fn pop_style() {
	sgl.pop_pipeline()

	mut ctx := context()
	if unsafe { ctx.cc == nil } {
		if ctx.cc.style_history.len() > 0 {
			style := ctx.cc.style_history.pop() or { panic(err) }
			set_style(style, mut ctx.cc)
		}
	}
}
module cc
// import gg
import sokol.sgl

pub fn push_matrix() {
	sgl.push_matrix()
}

pub fn pop_matrix() {
	sgl.pop_matrix()
}